


module riscv_bus_arbiter
    #(
        parameter DEVICE_1 = 1
    )
    (
        // *** SYSTEM PINS
        input CLK, input NRST,

        // *** IO
		

        // ***

    );