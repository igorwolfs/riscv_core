module core_cmem (
)


endmodule
