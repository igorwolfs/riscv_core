//! *************** PERIPHERAL CONFIGURATION ******************

`define INTERNAL_MEMORY	1